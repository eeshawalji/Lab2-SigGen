module sinegen #(
    parameter A_WIDTH = 8,
              D_WIDTH = 8
)(
    //interface signals
    input logic         clk,
    input logic         rst,
    input logic         en,
    input logic [D_WIDTH-1:0] incr,
    output logic [D_WIDTH-1:0] dout1,
    output logic [D_WIDTH-1:0] dout2
);

  logic [A_WIDTH-1:0] addr1;

counter addrCounter (
    .clk (clk),
    .rst (rst),
    .en (en),
    //.incr (incr),
    .count (addr1)
);

rom sineRom (
    .clk (clk),
    .addr1 (addr1),
    .dout1 (dout1),
    .addr2 (addr1+incr),
    .dout2 (dout2)
);


endmodule
